`include "components/uvm/comp_decomp_env.sv"

class comp_decomp_test extends uvm_test;
    
    `uvm_component_utils(comp_decomp_test)

    comp_decomp_env env;


    function new (string name = "comp_decomp_test", uvm_component parent=null);
        super.new(name,parent);
    endfunction

    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        env = comp_decomp_env::type_id::create("env", this);
    endfunction : build_phase

    virtual function void end_of_elaboration_phase(uvm_phase phase);
        print();
    endfunction

    function void report_phase(uvm_phase phase);
        uvm_report_server svr;

        super.report_phase(phase);

        svr = uvm_report_server::get_server();

        if (svr.get_severity_count(UVM_FATAL) + svr.get_severity_count(UVM_ERROR) > 0) begin
            `uvm_info(get_type_name(), "---------------------------------------", UVM_NONE)
            `uvm_info(get_type_name(), "----            TEST FAIL          ----", UVM_NONE)
            `uvm_info(get_type_name(), "---------------------------------------", UVM_NONE)
        end else begin   
            `uvm_info(get_type_name(), "---------------------------------------", UVM_NONE)
            `uvm_info(get_type_name(), "----           TEST PASS           ----", UVM_NONE)
            `uvm_info(get_type_name(), "---------------------------------------", UVM_NONE)
        end
    endfunction

endclass //comp_decomp_env extends uvm_tests